entity Adder_16b is
    port(
        a, b : in BIT_VECTOR(15 downto 0);
        cin  : in bit;
        s    : out BIT_VECTOR(15 downto 0);
        cout : out bit
    );
end Adder_16b;

architecture behav of Adder_16b is

begin

end architecture behav;
