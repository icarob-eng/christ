entity Reg_1b is -- D flip-flop
    port(
        input, write_en, clk : in  bit;
        output               : out bit
    );
end Reg_1b;


architecture behav of Reg_1b is

begin

end architecture behav;
