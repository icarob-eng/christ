entity Mux2x1_5b is
    port(
        i0, i1 : in  BIT_VECTOR(4 downto 0);
        s      : in  bit;
        o      : out BIT_VECTOR(4 downto 0)
    );
end Mux2x1_5b;


architecture behav of Mux2x1_5b is

begin

end architecture behav;
