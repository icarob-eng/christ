entity Mux2x1_3b is
    port(
        i0, i1 : in  BIT_VECTOR(2 downto 0);
        s      : in  bit;
        o      : out BIT_VECTOR(2 downto 0)
    );
end Mux2x1_3b;


architecture behav of Mux2x1_3b is

begin

end architecture behav;
